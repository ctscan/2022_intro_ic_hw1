module q3 (out, inp, clk);
  output reg out;
  input wire inp;
  input wire clk;
  
